* D:\Semester\FALL2021\CSE250\Lab2\20101065_Tanjim_Lab02\File2\20101065_TanjimReza_Lab2_File2.sch

* Schematics Version 9.2
* Thu Nov 04 01:32:31 2021



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "20101065_TanjimReza_Lab2_File2.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
