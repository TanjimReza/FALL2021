* C:\Users\Tanjim\Desktop\Lab3\Submission\20101065_TanjimRezaLab03File1.sch

* Schematics Version 9.2
* Sun Nov 14 22:02:06 2021



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "20101065_TanjimRezaLab03File1.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
